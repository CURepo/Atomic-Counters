/* *********************************
************************************
******* Atomic counter design ******
************************************
********************************* */


